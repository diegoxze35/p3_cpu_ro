LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
PACKAGE program IS
  CONSTANT EQ1_ADDR : INTEGER := 4;
  CONSTANT EQ2_ADDR : INTEGER := 25;
  CONSTANT EQ3_ADDR : INTEGER := 48;
END PACKAGE program;