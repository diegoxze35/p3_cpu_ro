LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY COMPARATOR_1_BIT IS
  PORT (
    A, B : IN STD_LOGIC;
    Gin, Ein, Lin : IN STD_LOGIC;
    Gout, Eout, Lout : OUT STD_LOGIC
  );
END COMPARATOR_1_BIT;
ARCHITECTURE Structural OF COMPARATOR_1_BIT IS
BEGIN
  Gout <= (A AND NOT B) OR ((A XNOR B) AND Gin);
  Eout <= (A XNOR B) AND Ein;
  Lout <= (NOT A AND B) OR ((A XNOR B) AND Lin);
END Structural;